//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Tue Jun 18 15:40:31 2024

module blk_mem_gen_3 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [10:0] ada;
input [7:0] dina;
input [10:0] adb;
input [7:0] dinb;

wire [7:0] dpb_inst_0_douta_w;
wire [7:0] dpb_inst_0_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[7:0],douta[7:0]}),
    .DOB({dpb_inst_0_doutb_w[7:0],doutb[7:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:0]}),
    .ADB({adb[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b1;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 8;
defparam dpb_inst_0.BIT_WIDTH_1 = 8;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h003C407E423C08040008080808080808007C12107C10120C0000000000000000;
defparam dpb_inst_0.INIT_RAM_01 = 256'h001C2222221C0014000002027E00000000223E2214081408003C424242420024;
defparam dpb_inst_0.INIT_RAM_02 = 256'h0000000000020408002222322C004C32003A464242420810005C22322A26221D;
defparam dpb_inst_0.INIT_RAM_03 = 256'h00223E2214084C3200223E22140800140044487844447A3E003A443C04380038;
defparam dpb_inst_0.INIT_RAM_04 = 256'h003C42423C004C32004834322A261609001C2222221C14000022262A32224C32;
defparam dpb_inst_0.INIT_RAM_05 = 256'h001C2A281C0A2A1C0018242418004C32003A464242420024007C22223C22223C;
defparam dpb_inst_0.INIT_RAM_06 = 256'h003C023E427C403C003A443C04380010003A443C04381020003A443C04380028;
defparam dpb_inst_0.INIT_RAM_07 = 256'h000000004C32000010081C222020221C0026243C26241E08003E203E203E0804;
defparam dpb_inst_0.INIT_RAM_08 = 256'h0024247E247E2424000000000024242400080008080808080000000000000000;
defparam dpb_inst_0.INIT_RAM_09 = 256'h0000000000100804003A444A30484830004626100864620000083C0A1C281E08;
defparam dpb_inst_0.INIT_RAM_0A = 256'h000008083E08080000082A1C3E1C2A0800201008080810200004081010100804;
defparam dpb_inst_0.INIT_RAM_0B = 256'h00402010080402000008000000000000000000007E0000001008080000000000;
defparam dpb_inst_0.INIT_RAM_0C = 256'h003C42021C02423C007E40300C02423C003E080808281808003C42625A46423C;
defparam dpb_inst_0.INIT_RAM_0D = 256'h001010100804427E003C42427C40201C003844020478407E0004047E24140C04;
defparam dpb_inst_0.INIT_RAM_0E = 256'h10080800000800000000080000080000003804023E42423C003C42423C42423C;
defparam dpb_inst_0.INIT_RAM_0F = 256'h001000100C02423C006030180C1830600000007E007E000000060C1830180C06;
defparam dpb_inst_0.INIT_RAM_10 = 256'h001C22404040221C007C22223C22227C004242427E422418001E204C564A221C;
defparam dpb_inst_0.INIT_RAM_11 = 256'h001C22424E40221C004040407840407E007E40407840407E0078242222222478;
defparam dpb_inst_0.INIT_RAM_12 = 256'h0042444870484442003844040404040E001C08080808081C004242427E424242;
defparam dpb_inst_0.INIT_RAM_13 = 256'h003C42424242423C004242464A526242004242425A5A6642007E404040404040;
defparam dpb_inst_0.INIT_RAM_14 = 256'h003C42023C40423C004244487C42427C003A444A4242423C004040407C42427C;
defparam dpb_inst_0.INIT_RAM_15 = 256'h0042665A5A4242420018182424424242003C424242424242000808080808083E;
defparam dpb_inst_0.INIT_RAM_16 = 256'h003C20202020203C007E40201804027E000808081C2222220042422418244242;
defparam dpb_inst_0.INIT_RAM_17 = 256'hFF000000000000000000000000221408003C04040404043C0002040810204000;
defparam dpb_inst_0.INIT_RAM_18 = 256'h003C4240423C0000005C6242625C4040003A443C043800000000000000040810;
defparam dpb_inst_0.INIT_RAM_19 = 256'h3C023A46463A0000001010107C10120C003C407E423C0000003A4642463A0202;
defparam dpb_inst_0.INIT_RAM_1A = 256'h004468504844404038440404040C0004001C08080818000800424242625C4040;
defparam dpb_inst_0.INIT_RAM_1B = 256'h003C4242423C000000424242625C00000049494949760000001C080808080818;
defparam dpb_inst_0.INIT_RAM_1C = 256'h007C023C403E000000404040625C000002023A46463A000040405C62625C0000;
defparam dpb_inst_0.INIT_RAM_1D = 256'h00364949494100000018244242420000003A464242420000000C1210107C1010;
defparam dpb_inst_0.INIT_RAM_1E = 256'h000C10102010100C007E2018047E00003C023A46424200000042241824420000;
defparam dpb_inst_0.INIT_RAM_1F = 256'h003E0008083E0808000000000006493000300808040808300008080800080808;
defparam dpb_inst_0.INIT_RAM_20 = 256'h1C086B7F6B081C1C00081C3E7F3E1C0800081C3E7F7F360008083E7F7F3E1C08;
defparam dpb_inst_0.INIT_RAM_21 = 256'h3C201008040810203C040810201008043C42A59981A5423C3C4299A581A5423C;
defparam dpb_inst_0.INIT_RAM_22 = 256'h000C120A0C10120C003030101814126140203C22223C223C0000394646390000;
defparam dpb_inst_0.INIT_RAM_23 = 256'h000814223E221408000202021212522C000C021C10080616000608103E100806;
defparam dpb_inst_0.INIT_RAM_24 = 256'h0020203A24242424004224181010102000444A5060504840001C222220202000;
defparam dpb_inst_0.INIT_RAM_25 = 256'h00141414543E000000182442422418000C021C2018201C080010181412320000;
defparam dpb_inst_0.INIT_RAM_26 = 256'h001824242464020008080808483E000000003048483E00000020203824241800;
defparam dpb_inst_0.INIT_RAM_27 = 256'h0036494941220000000808081C2A2A49002314081462000000081C2A2A2A1C08;
defparam dpb_inst_0.INIT_RAM_28 = 256'h007E20100C10207E000008003E000800001030501010101E006322634141221C;
defparam dpb_inst_0.INIT_RAM_29 = 256'h0040207F087F0201201008081010080400007F221408000000004C32004C3200;
defparam dpb_inst_0.INIT_RAM_2A = 256'h00003649493600006322227F4141221C004225120824523F000408103E040810;
defparam dpb_inst_0.INIT_RAM_2B = 256'h3C429DA1A19D423C0022552A142A5522003C021C221C201E0040605048040200;
defparam dpb_inst_0.INIT_RAM_2C = 256'h3C66A9B9A5A57A3C00081C2A282A1C080A0A0A0A3A4A4A3E0042241824182442;
defparam dpb_inst_0.INIT_RAM_2D = 256'h004B444A784444780000000000FC02FCF804FC02FC0304FF5F607B646263605F;
defparam dpb_inst_0.INIT_RAM_2E = 256'h000000000E08080E081C081C2222221C00609090700A060E8649291668848261;
defparam dpb_inst_0.INIT_RAM_2F = 256'h22362A2222221408143E142A1C0814082214082A1C081408FFF7FFF7F3DDE3FF;
defparam dpb_inst_0.INIT_RAM_30 = 256'h001C040404000000000000001010101C002050200000000000083E083E081422;
defparam dpb_inst_0.INIT_RAM_31 = 256'h0010080C023E0000000804027E027E0000000018180000000010200000000000;
defparam dpb_inst_0.INIT_RAM_32 = 256'h0024140C3E040000003E08083E000000000804223E0800000004140C04020000;
defparam dpb_inst_0.INIT_RAM_33 = 256'h000C022A2A000000003C041C043C0000003E04041C000000001014123E100000;
defparam dpb_inst_0.INIT_RAM_34 = 256'h0008040202427E1000084828180804020020101816027E00000000003E000000;
defparam dpb_inst_0.INIT_RAM_35 = 256'h000808087F087F080044221212127E1000044424140C7E04003E080808083E00;
defparam dpb_inst_0.INIT_RAM_36 = 256'h0010080424247E24007E020202027E000010080808483E200010080442223E20;
defparam dpb_inst_0.INIT_RAM_37 = 256'h0010080402224200000E101012117E100022140804023E000038040262026000;
defparam dpb_inst_0.INIT_RAM_38 = 256'h001008087E003C000008040252525200001008087E0838040010080C52223E20;
defparam dpb_inst_0.INIT_RAM_39 = 256'h0022140814023E00007E000000003C0000100808087E08080010121418101010;
defparam dpb_inst_0.INIT_RAM_3A = 256'h003E4040407E4040004242424408100000201008080808080050321408047E10;
defparam dpb_inst_0.INIT_RAM_3B = 256'h000408182402027E0008494908087F080001010244281000001804020202027E;
defparam dpb_inst_0.INIT_RAM_3C = 256'h000E10107E107E00004020140814020200027E424020100800027C003C003C40;
defparam dpb_inst_0.INIT_RAM_3D = 256'h00080402027E003C003E02023E02023E007F040404043C0000101014127E1010;
defparam dpb_inst_0.INIT_RAM_3E = 256'h007E424242427E00006050484440404000585452505050100010080444444444;
defparam dpb_inst_0.INIT_RAM_3F = 256'h0000000000205020000000000020481000780402020060000008040242427E00;

endmodule //blk_mem_gen_3
